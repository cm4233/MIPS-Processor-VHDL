--VHDL Code for the ALU (Arithmetic and Logic Unit) of the MIPS Processor--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity alu is
---------//ports//---------
PORT (
SrcA: in STD_LOGIC_VECTOR(31 DOWNTO 0);
SrcB: in STD_LOGIC_VECTOR(31 DOWNTO 0);
ALUControl: in STD_LOGIC_VECTOR(2 DOWNTO 0);

Zero: out STD_LOGIC;
GreatThan: out STD_LOGIC;
LessThan: out STD_LOGIC;
ALUResult: out STD_LOGIC_VECTOR(31 DOWNTO 0));
--------------------------
end alu;

architecture Behavioral of alu is
------//signals//-------------
signal z: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal shiftleft: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal shiftright: STD_LOGIC_VECTOR(31 DOWNTO 0);
----------------------------
begin
----------//code//---------
z<=SrcA-SrcB;
--leftshift--
WITH SrcB(15 DOWNTO 0) SELECT
    shiftleft<=	SrcA(30 DOWNTO 0) & '0' WHEN "0000000000000001",
	SrcA(29 DOWNTO 0) & "00" WHEN "0000000000000010",
	SrcA(28 DOWNTO 0) & "000" WHEN "0000000000000011",
	SrcA(27 DOWNTO 0) & "0000" WHEN "0000000000000100",
	SrcA(26 DOWNTO 0) & "00000" WHEN "0000000000000101",
	SrcA(25 DOWNTO 0) & "000000" WHEN "0000000000000110",
	SrcA(24 DOWNTO 0) & "0000000" WHEN "0000000000000111",
	SrcA(23 DOWNTO 0) & "00000000" WHEN "0000000000001000",
	SrcA(22 DOWNTO 0) & "000000000" WHEN "0000000000001001",
	SrcA(21 DOWNTO 0) & "0000000000" WHEN "0000000000001010",
	SrcA(20 DOWNTO 0) & "00000000000" WHEN "0000000000001011",
	SrcA(19 DOWNTO 0) & "000000000000" WHEN "0000000000001100",
	SrcA(18 DOWNTO 0) & "0000000000000" WHEN "0000000000001101",
	SrcA(17 DOWNTO 0) & "00000000000000" WHEN "0000000000001110",
	SrcA(16 DOWNTO 0) & "000000000000000" WHEN "0000000000001111",
	SrcA(15 DOWNTO 0) & "0000000000000000" WHEN "0000000000010000",
	SrcA(14 DOWNTO 0) & "00000000000000000" WHEN "0000000000010001",
	SrcA(13 DOWNTO 0) & "000000000000000000" WHEN "0000000000010010",
	SrcA(12 DOWNTO 0) & "0000000000000000000" WHEN "0000000000010011",
	SrcA(11 DOWNTO 0) & "00000000000000000000" WHEN "0000000000010100",
	SrcA(10 DOWNTO 0) & "000000000000000000000" WHEN "0000000000010101",
	SrcA(9 DOWNTO 0) &  "0000000000000000000000" WHEN "0000000000010110",
	SrcA(8 DOWNTO 0) &  "00000000000000000000000" WHEN "0000000000010111",
	SrcA(7 DOWNTO 0) &  "000000000000000000000000" WHEN "0000000000011000",
	SrcA(6 DOWNTO 0) &  "0000000000000000000000000" WHEN "0000000000011001",
	SrcA(5 DOWNTO 0) &  "00000000000000000000000000" WHEN "0000000000011010",
	SrcA(4 DOWNTO 0) &  "000000000000000000000000000" WHEN "0000000000011011",
	SrcA(3 DOWNTO 0) &  "0000000000000000000000000000" WHEN "0000000000011100",
	SrcA(2 DOWNTO 0) &  "00000000000000000000000000000" WHEN "0000000000011101",
	SrcA(1 DOWNTO 0) &  "000000000000000000000000000000" WHEN "0000000000011110",
	SrcA(0) &           "0000000000000000000000000000000" WHEN "0000000000011111",
	SrcA WHEN OTHERS;
--rightshift--
WITH SrcB(15 DOWNTO 0) SELECT
    shiftright<=	'0' & SrcA(31 DOWNTO 1)  WHEN "0000000000000001",
	"00" & SrcA(31 DOWNTO 2)   WHEN "0000000000000010",
	"000" & SrcA(31 DOWNTO 3)   WHEN "0000000000000011",
	"0000" & SrcA(31 DOWNTO 4)   WHEN "0000000000000100",
	"00000" & SrcA(31 DOWNTO 5)   WHEN "0000000000000101",
	"000000" & SrcA(31 DOWNTO 6)   WHEN "0000000000000110",
	"0000000" & SrcA(31 DOWNTO 7)   WHEN "0000000000000111",
	"00000000" & SrcA(31 DOWNTO 8)   WHEN "0000000000001000",
	"000000000" & SrcA(31 DOWNTO 9)   WHEN "0000000000001001",
	"0000000000" & SrcA(31 DOWNTO 10)   WHEN "0000000000001010",
	"00000000000" & SrcA(31 DOWNTO 11)   WHEN "0000000000001011",
	"000000000000" & SrcA(31 DOWNTO 12)   WHEN "0000000000001100",
	"0000000000000" & SrcA(31 DOWNTO 13)   WHEN "0000000000001101",
	"00000000000000" & SrcA(31 DOWNTO 14)   WHEN "0000000000001110",
	"000000000000000" & SrcA(31 DOWNTO 15)   WHEN "0000000000001111",
	"0000000000000000" & SrcA(31 DOWNTO 16)   WHEN "0000000000010000",
	"00000000000000000" & SrcA(31 DOWNTO 17)   WHEN "0000000000010001",
	"000000000000000000" & SrcA(31 DOWNTO 18)   WHEN "0000000000010010",
	"0000000000000000000" & SrcA(31 DOWNTO 19)   WHEN "0000000000010011",
	"00000000000000000000" & SrcA(31 DOWNTO 20)   WHEN "0000000000010100",
	"000000000000000000000" & SrcA(31 DOWNTO 21)   WHEN "0000000000010101",
	"0000000000000000000000" & SrcA(31 DOWNTO 22)    WHEN "0000000000010110",
	"00000000000000000000000" & SrcA(31 DOWNTO 23)    WHEN "0000000000010111",
	"000000000000000000000000" & SrcA(31 DOWNTO 24)    WHEN "0000000000011000",
	"0000000000000000000000000" & SrcA(31 DOWNTO 25)    WHEN "0000000000011001",
	"00000000000000000000000000" & SrcA(31 DOWNTO 26)    WHEN "0000000000011010",
	"000000000000000000000000000" & SrcA(31 DOWNTO 27)    WHEN "0000000000011011",
	"0000000000000000000000000000" & SrcA(31 DOWNTO 28)    WHEN "0000000000011100",
	"00000000000000000000000000000" & SrcA(31 DOWNTO 29)    WHEN "0000000000011101",
	"000000000000000000000000000000" & SrcA(31 DOWNTO 30)    WHEN "0000000000011110",
	"0000000000000000000000000000000" & SrcA(31)             WHEN "0000000000011111",
	SrcA WHEN OTHERS;
-------------------------------------
with ALUControl select
ALUResult <= 	SrcA+SrcB when "000",
					SrcA-SrcB when "001",
					SrcA and SrcB when "010",
					SrcA or SrcB when "011",
					SrcA nor SrcB when "100",
					shiftleft when "101",
					shiftright when "110",
					SrcA+SrcB when others;	

with z select
Zero <= 	'1' when x"00000000",
			'0' when others;	
with z(31) select
LessThan <= 	'1' when '1',
					'0' when others;
with z select					
GreatThan <= 	'0' when x"00000000",
					--not z(31) when others;
					'1' when others;
----------------------------
end Behavioral;

