--VHDL Code for the IM (Instruction Memory) of the MIPS Processor--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity instructionmemory is
---------//ports//--------------------------------------
PORT (address: in STD_LOGIC_VECTOR(31 DOWNTO 0);
 	   data: out STD_LOGIC_VECTOR(31 DOWNTO 0));
-----------------------------------------------
end instructionmemory;

architecture Behavioral of instructionmemory is
--------//signals//------------------------
TYPE rom IS ARRAY (0 TO 220) OF STD_LOGIC_VECTOR(31 DOWNTO 0); 
CONSTANT imem: 
rom:=rom'(
---------Instruction memory loaded with RC5 encrytion and decryption code------
-----------ENCRYPT SKEY GEN-----------------------------
-------------UKEY FROM MEM---------------
"00011100000110010000000000100010",--LW R25,34(R0) i0
"00100000000110010000000000011100",--SW R25,28(R0)
"00011100000110010000000000100011",--LW R25,35(R0)
"00100000000110010000000000011101",--SW R25,29(R0)
"00011100000110010000000000100100",--LW R25,36(R0)
"00100000000110010000000000011110",--SW R25,30(R0)
"00011100000110010000000000100101",--LW R25,37(R0)
"00100000000110010000000000011111",--SW R25,31(R0) i7
-----------------------------------------
"00000100000110000000000001001110", --	ADDI R24,R0,#4E h i8
"00000100000101100000000000011010", --	ADDI R22,R0,#1A h
"00000100000101110000000000000100", --	ADDI R23,R0,#04 h 
"00000100000100110000000000100000", --	ADDI R19,R0,#20 h
"00000000000000000010100000010000", -- ADD R5,R0,R0
"00000000000000000010000000010000", -- ADD R4,R0,R0
"00000000000000000000100000010000", -- ADD R1,R0,R0
"00011100010001100000000000000000", --LW R6,0(R2)  LOOP
"00000000100001010011100000010000", -- ADD R7 R4 R5
"00000000111001100100000000010000", -- ADD R8 R7 R6
"00010101000010010000000000000011", --SHL R9 R8 3
"00011001000010100000000000011101", --SHR R10 R8 1D hex
"00000001001010100101100000010011", --OR R11 R9 R10
"00100000010010110000000000000000", --SW R11 ,0(R2)
"00000000000010110010000000010000", -- ADD R4 R11 R0
"00000000101010110110000000010000", -- ADD R12 R11 R5
"00011100011011010000000000011100", --LW R13 ,28(R3)
"00000001100011010111000000010000", -- ADD R14 R13 R12
"00001101100011110000000000011111", --ANDI R15,R12,#1Fh
"00000000000000001000000000010000",	--ADD R16,R0,R0
"00000000000011101000100000010000",	--ADD R17,R14,R0
"00101000000011110000000000001010",	--BEQ R15,R0,10
"00000000000011101000000000010000", --ADD R16,R14,R0
"00000000000011101000100000010000",	--ADD R17,R14,R0
"00000000000011111001000000010000", --ADD R18,R15,R0 //r9=r15,r10=r18
"00010110000100000000000000000001", --SHL R16,R16,#1h //r11=r16
"00001010010100100000000000000001", --SUBI R18,R18,#1h
"00101100000100101111111111111101", --BNE R18,R0,#(-3)
"00000010011011111010000000010001", --SUB R20,R19,R15 //r13=r20 r12=r19//LOAD R19 20hex
"00011010001100010000000000000001", --SHR R17,R17,#1h //r14=r17
"00001010100101000000000000000001", --SUBI R20,R20,1
"00101100000101001111111111111101", --BNE R20 ,R0, -3
"00000010000100011010100000010011", --OR R21 R17 R16
"00000000000101010010100000010000", -- ADD R5 R0 R21
"00100000011101010000000000011100", --SW R21 ,28(R3)
"00000100011000110000000000000001", --ADDI R3 R3 1
"00101100011101110000000000000001", --BNE R3,R23,1
"00000000000000000001100000010000", -- ADD R3,R0,R0 
"00000100010000100000000000000001", --ADDI R2 R2 1
"00101100010101100000000000000001", --BNE R2 R22,1
"00000000000000000001000000010000", -- ADD R2,R0,R0 
"00000100001000010000000000000001", --ADDI R1 R1 1
"00101100001110001111111111011100", --BNE R1 R24,-36 LOOP
"00101000000000000000000000000000", --BEQ R0 R0 0 i51
-----------END OF ENCRYPT SKEY GEN----------
-------encryption----
"00011100000110100000000000000000",	--LW R26,0(R0) i52
"00011100000110110000000000000001", --LW R27,1(R0)
"00011100000000010000000000100000", --LW R1,32(R0)
"00011100000000100000000000100001", --LW R2,33(R0)
"00000000001110100000100000010000", --ADD R1,R1,R26 
"00000000010110110001000000010000", --ADD R2,R2,R27 
"00000100000000110000000000000001", --ADDI R3,R0,#1h
"00000100000011000000000000100000", --ADDI R12,R0,#20h
"00000100000101010000000000001101", --ADDI R21,R0,#Dh
"00000000010000100010000000010100", --NOR R4,R2,R2
"00000000001000010010100000010100", --NOR R5,R1,R1
"00000000100000010011000000010010", --AND R6,R1,R4
"00000000010001010011100000010010", --AND R7,R5,R2
"00000000111001100100000000010011", --OR R8,R6,R7
"00001100010010010000000000011111", --ANDI R9,R2,#1Fh i66
------------------------------------------------------42down
"00000000000000000111000000010000",	--ADD R14,R0,R0 i67
"00000000000010000101100000010000",	--ADD R11,R8,R0
"00101000000010010000000000001010",	--BEQ R9,R0,10
"00000000000010000101100000010000", --ADD R11,R8,R0
"00000000000010000111000000010000",	--ADD R14,R8,R0 i71
------------------------------------------------------37down
"00000000000010010101000000010000", --ADD R10,R9,R0 i72
"00010101011010110000000000000001", --SHL R11,R11,#1h
"00001001010010100000000000000001", --SUBI R10,R10,#1h
"00101100000010101111111111111101", --BNE R10,R0,#(-3)
"00000001100010010110100000010001", --SUB R13,R12,R9
"00011001110011100000000000000001", --SHR R14,R14,#1h
"00001001101011010000000000000001", --SUBI R13,R13,1
"00101100000011011111111111111101", --BNE R13 ,R0, -3
"00000001011011100111100000010011", --OR R15 R14 R11
"00010100011100000000000000000001", --SHL R16 R3 1
"00000110000100010000000000000001", --ADDI R17 R16 1
"00011110000100110000000000000000", --LW R19 0(R16)
"00000010011011110000100000010000", --ADD R1 R15 R19
"00000000010000100010000000010100", --NOR R4,R2,R2
"00000000001000010010100000010100", --NOR R5,R1,R1
"00000000100000010011000000010010", --AND R6,R1,R4
"00000000010001010011100000010010", --AND R7,R5,R2
"00000000111001100100000000010011", --OR R8,R6,R7
"00001100001010010000000000011111",  --ANDI R9,R1,#1Fh i90
------------------------------------------------------18down
"00000000000000000111000000010000",	--ADD R14,R0,R0 i91
"00000000000010000101100000010000",	--ADD R11,R8,R0
"00101000000010010000000000001010",	--BEQ R9,R0,10
"00000000000010000101100000010000", --ADD R11,R8,R0
"00000000000010000111000000010000",	--ADD R14,R8,R0 i95
------------------------------------------------------
"00000000000010010101000000010000", --ADD R10,R9,R0 i96
"00010101011010110000000000000001", --SHL R11,R11,#1h
"00001001010010100000000000000001",  --SUBI R10,R10,#1h
"00101100000010101111111111111101", --BNE R10,R0,#(-3)
"00000001100010010110100000010001", --SUB R13,R12,R9
"00011001110011100000000000000001", --SHR R14,R14,#1h
"00001001101011010000000000000001", --SUBI R13,R13,1
"00101100000011011111111111111101", --BNE R13 ,R0, -3
"00000001011011100111100000010011", --OR R15 R14 R11
"00011110001101000000000000000000", --LW R20 0(R17)
"00000010100011110001000000010000", --ADD R2 R15 R20
"00000100011000110000000000000001", --ADDI R3 R3 1
"00101110101000111111111111010000", --BNE R3 R21 (-48)
"00101000000000001111111111111111", --BEQ R0 R0 -1 infinite loop i109
-----------------end of encryption-----------------------------------------
-----------DECRYPT SKEY GEN-----------------------------
-------------UKEY FROM MEM---------------
"00011100000110010000000000100010",--LW R25,34(R0) i110
"00100000000110010000000000011100",--SW R25,28(R0)
"00011100000110010000000000100011",--LW R25,35(R0)
"00100000000110010000000000011101",--SW R25,29(R0)
"00011100000110010000000000100100",--LW R25,36(R0)
"00100000000110010000000000011110",--SW R25,30(R0)
"00011100000110010000000000100101",--LW R25,37(R0)
"00100000000110010000000000011111",--SW R25,31(R0)
-----------------------------------------
"00000100000110000000000001001110", --	ADDI R24,R0,#4E h
"00000100000101100000000000011010", --	ADDI R22,R0,#1A h
"00000100000101110000000000000100", --	ADDI R23,R0,#04 h 
"00000100000100110000000000100000", --	ADDI R19,R0,#20 h
"00000000000000000010100000010000", -- ADD R5,R0,R0
"00000000000000000010000000010000", -- ADD R4,R0,R0
"00000000000000000000100000010000", -- ADD R1,R0,R0
"00011100010001100000000000000000", --LW R6,0(R2)  LOOP
"00000000100001010011100000010000", -- ADD R7 R4 R5
"00000000111001100100000000010000", -- ADD R8 R7 R6
"00010101000010010000000000000011", --SHL R9 R8 3
"00011001000010100000000000011101", --SHR R10 R8 1D hex
"00000001001010100101100000010011", --OR R11 R9 R10
"00100000010010110000000000000000", --SW R11 ,0(R2)
"00000000000010110010000000010000", -- ADD R4 R11 R0
"00000000101010110110000000010000", -- ADD R12 R11 R5
"00011100011011010000000000011100", --LW R13 ,28(R3)
"00000001100011010111000000010000", -- ADD R14 R13 R12
"00001101100011110000000000011111", --ANDI R15,R12,#1Fh
"00000000000000001000000000010000",	--ADD R16,R0,R0
"00000000000011101000100000010000",	--ADD R17,R14,R0
"00101000000011110000000000001010",	--BEQ R15,R0,10
"00000000000011101000000000010000", --ADD R16,R14,R0
"00000000000011101000100000010000",	--ADD R17,R14,R0
"00000000000011111001000000010000", --ADD R18,R15,R0 //r9=r15,r10=r18
"00010110000100000000000000000001", --SHL R16,R16,#1h //r11=r16
"00001010010100100000000000000001", --SUBI R18,R18,#1h
"00101100000100101111111111111101", --BNE R18,R0,#(-3)
"00000010011011111010000000010001", --SUB R20,R19,R15 //r13=r20 r12=r19//LOAD R19 20hex
"00011010001100010000000000000001", --SHR R17,R17,#1h //r14=r17
"00001010100101000000000000000001", --SUBI R20,R20,1
"00101100000101001111111111111101", --BNE R20 ,R0, -3
"00000010000100011010100000010011", --OR R21 R17 R16
"00000000000101010010100000010000", -- ADD R5 R0 R21
"00100000011101010000000000011100", --SW R21 ,28(R3)
"00000100011000110000000000000001", --ADDI R3 R3 1
"00101100011101110000000000000001", --BNE R3,R23,1
"00000000000000000001100000010000", -- ADD R3,R0,R0 
"00000100010000100000000000000001", --ADDI R2 R2 1
"00101100010101100000000000000001", --BNE R2 R22,1
"00000000000000000001000000010000", -- ADD R2,R0,R0 
"00000100001000010000000000000001", --ADDI R1 R1 1
"00101100001110001111111111011100", --BNE R1 R24,-36 LOOP
"00101000000000000000000000000000", --BEQ R0 R0 0
-----------END OF DECRYPT SKEY GEN----------
-------decryption-----------------------------
"00011100000000010000000000100000", --LWR1,32(R0)
"00011100000000100000000000100001", --LWR2 33(R0)
"00000100000000110000000000001101", --ADDI R3 R0 #DH
"00000100000001000000000000000001", --ADDI R4 R0 #1H
"00000100000001010000000000100000", --ADDI R5 R0 #20H
"00010100011001100000000000000001", --SHL R6 R3 #1H --
"00001000110001110000000000000001", --SUBI R7 R6 #1H
"00001000110010000000000000000010", --SUBI R8 R6 #2H
"00011100111010010000000000000000", --LWR9 0(R7)
"00011101000010100000000000000000", --LWR10,0(R8)
"00000000010010010101100000010001", --SUB R11 R2 R9 
"00001100001011000000000000011111", --ANDI R12 R1 #1FH
"00000001100000000110100000010000", --ADD R13 R12 R0
"00000001011000000111000000010000", --ADD R14 R11 R0
"00000000000000001000000000010000", --ADD R16 R0 R0
"00101000000011000000000000001000", --BEQ R12 R0 8
"00000001011000000111000000010000", --ADD R14 R11 R0
"00000001011000001000000000010000", --ADD R16 R11 R0
"00011001110011100000000000000001", --SHR R14 R14 1
"00001001101011010000000000000001", --SUBI R13 R13 1
"00101100000011011111111111111101", --BNE R13 R0 -3
"00000000101011000111100000010001", --SUB R15 R5 R12
"00010110000100000000000000000001", --SHL R16 R16 1
"00001001111011110000000000000001", --SUBI R15 R15 1
"00101100000011111111111111111101", --BNE R15 R0 -3
"00000010000011101000100000010011", --OR R17 R16 R14
"00000010001100011001000000010100", --NOR R18 R17 R17
"00000000001000011001100000010100", --NOR R19 R1 R1
"00000000001100101010000000010010", --AND R20 R1 R18
"00000010001100111010100000010010", --AND R21 R17 R19
"00000010100101010001000000010011", --OR R2 R20 R21
"00000000001010100101100000010001", --SUB R11 R1 R10
"00001100010011000000000000011111", --ANDI R12 R2 #1FH
"00000001100000000110100000010000", --ADD R13 R12 R0
"00000001011000000111000000010000", --ADD R14 R11 R0
"00000000000000001000000000010000", --ADD R16 R0 R0
"00101000000011000000000000001000", --BEQ R12 R0 8
"00000001011000000111000000010000", --ADD R14 R11 R0
"00000001011000001000000000010000", --ADD R16 R11 R0
"00011001110011100000000000000001", --SHR R14 R14 1
"00001001101011010000000000000001", --SUBI R13 R13 1
"00101100000011011111111111111101", --BNE R13 R0 -3
"00000000101011000111100000010001", --SUB R15 R5 R12
"00010110000100000000000000000001", --SHL R16 R16 1
"00001001111011110000000000000001", --SUBI R15 R15 1
"00101100000011111111111111111101", --BNE R15 R0 -3
"00000010000011101000100000010011", --OR R17 R16 R14
"00000010001100011001000000010100", --NOR R18 R17 R17
"00000000010000101001100000010100", --NOR R19 R2 R2
"00000010011100011010000000010010", --AND R20 R19 R17
"00000000010100101010100000010010", --AND R21 R2 R18
"00000010100101010000100000010011", --OR R1 R20 R21
"00001000011000110000000000000001", --SUBI R3 R3 1
"00101100100000111111111111001111", --BNE R3 R4 -49
"00011100000000110000000000000000", --LWR3,0(R0)
"00000000001000110000100000010001", --SUB R1 R1 R3
"00011100000001000000000000000001", --LWR4 1(R0)
"00000000010001000001000000010001", --SUB R2 R2 R4
"00101000000000001111111111111111"); --BEQ R0 R0 -1 infinite loop
-------end of decryption----------------------
--------------------------------------
begin
---------//code//-------------------
data<=imem(CONV_INTEGER(address));
------------------------------------
end Behavioral;

