--VHDL Code for the ALU (Arithmetic and Logic Unit) of the MIPS Processor--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity alu is
---------//ports//---------
PORT (
SrcA: in STD_LOGIC_VECTOR(31 DOWNTO 0);--Operand 1
SrcB: in STD_LOGIC_VECTOR(31 DOWNTO 0);--Operand 2
ALUControl: in STD_LOGIC_VECTOR(2 DOWNTO 0);--The ALU operation to be performed on the operands. Controlled by CU.

Zero: out STD_LOGIC;--'1' if Operand 1 & 2 are equal. Used mainly for BEQ instruction
GreatThan: out STD_LOGIC;--'1' if Op1>Op2. Used for BGT instruction
LessThan: out STD_LOGIC;--'1' if Op1<Op2. Used for BLT instruction
ALUResult: out STD_LOGIC_VECTOR(31 DOWNTO 0));--The result of the ALU operation
--------------------------
end alu;

architecture Behavioral of alu is
------//intermediate signals//-------------
signal z: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal shiftleft: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal shiftright: STD_LOGIC_VECTOR(31 DOWNTO 0);
----------------------------
begin
----------//code//---------
z<=SrcA-SrcB;
--leftshift--
with SrcB select
	shiftleft<=	
	SrcA WHEN x"00000000",
	SrcA(30 DOWNTO 0) & '0' WHEN x"00000001",
	SrcA(29 DOWNTO 0) & "00" WHEN x"00000002",
	SrcA(28 DOWNTO 0) & "000" WHEN x"00000003",
	SrcA(27 DOWNTO 0) & "0000" WHEN x"00000004",
	SrcA(26 DOWNTO 0) & "00000" WHEN x"00000005",
	SrcA(25 DOWNTO 0) & "000000" WHEN x"00000006",
	SrcA(24 DOWNTO 0) & "0000000" WHEN x"00000007",
	SrcA(23 DOWNTO 0) & "00000000" WHEN x"00000008",
	SrcA(22 DOWNTO 0) & "000000000" WHEN x"00000009",
	SrcA(21 DOWNTO 0) & "0000000000" WHEN x"0000000A",
	SrcA(20 DOWNTO 0) & "00000000000" WHEN x"0000000B",
	SrcA(19 DOWNTO 0) & "000000000000" WHEN x"0000000C",
	SrcA(18 DOWNTO 0) & "0000000000000" WHEN x"0000000D",
	SrcA(17 DOWNTO 0) & "00000000000000" WHEN x"0000000E",
	SrcA(16 DOWNTO 0) & "000000000000000" WHEN x"0000000F",
	SrcA(15 DOWNTO 0) & "0000000000000000" WHEN x"00000010",
	SrcA(14 DOWNTO 0) & "00000000000000000" WHEN x"00000011",
	SrcA(13 DOWNTO 0) & "000000000000000000" WHEN x"00000012",
	SrcA(12 DOWNTO 0) & "0000000000000000000" WHEN x"00000013",
	SrcA(11 DOWNTO 0) & "00000000000000000000" WHEN x"00000014",
	SrcA(10 DOWNTO 0) & "000000000000000000000" WHEN x"00000015",
	SrcA(9 DOWNTO 0) &  "0000000000000000000000" WHEN x"00000016",
	SrcA(8 DOWNTO 0) &  "00000000000000000000000" WHEN x"00000017",
	SrcA(7 DOWNTO 0) &  "000000000000000000000000" WHEN x"00000018",
	SrcA(6 DOWNTO 0) &  "0000000000000000000000000" WHEN x"00000019",
	SrcA(5 DOWNTO 0) &  "00000000000000000000000000" WHEN x"0000001A",
	SrcA(4 DOWNTO 0) &  "000000000000000000000000000" WHEN x"0000001B",
	SrcA(3 DOWNTO 0) &  "0000000000000000000000000000" WHEN x"0000001C",
	SrcA(2 DOWNTO 0) &  "00000000000000000000000000000" WHEN x"0000001D",
	SrcA(1 DOWNTO 0) &  "000000000000000000000000000000" WHEN x"0000001E",
	SrcA(0) &           "0000000000000000000000000000000" WHEN x"0000001F",
	x"00000000" WHEN OTHERS;
--rightshift--
WITH SrcB SELECT
   shiftright<=
	SrcA WHEN x"00000000",
	'0' & SrcA(31 DOWNTO 1) WHEN x"00000001",
	"00" & SrcA(31 DOWNTO 2) WHEN x"00000002",
	"000" & SrcA(31 DOWNTO 3) WHEN x"00000003",
	"0000" & SrcA(31 DOWNTO 4) WHEN x"00000004",
	"00000" & SrcA(31 DOWNTO 5) WHEN x"00000005",
	"000000" & SrcA(31 DOWNTO 6) WHEN x"00000006",
	"0000000" & SrcA(31 DOWNTO 7) WHEN x"00000007",
	"00000000" & SrcA(31 DOWNTO 8) WHEN x"00000008",
	"000000000" & SrcA(31 DOWNTO 9) WHEN x"00000009",
	"0000000000" & SrcA(31 DOWNTO 10) WHEN x"0000000A",
	"00000000000" & SrcA(31 DOWNTO 11) WHEN x"0000000B",
	"000000000000" & SrcA(31 DOWNTO 12) WHEN x"0000000C",
	"0000000000000" & SrcA(31 DOWNTO 13) WHEN x"0000000D",
	"00000000000000" & SrcA(31 DOWNTO 14) WHEN x"0000000E",
	"000000000000000" & SrcA(31 DOWNTO 15) WHEN x"0000000F",
	"0000000000000000" & SrcA(31 DOWNTO 16) WHEN x"00000010",
	"00000000000000000" & SrcA(31 DOWNTO 17) WHEN x"00000011",
	"000000000000000000" & SrcA(31 DOWNTO 18) WHEN x"00000012",
	"0000000000000000000" & SrcA(31 DOWNTO 19) WHEN x"00000013",
	"00000000000000000000" & SrcA(31 DOWNTO 20) WHEN x"00000014",
	"000000000000000000000" & SrcA(31 DOWNTO 21) WHEN x"00000015",
	"0000000000000000000000" & SrcA(31 DOWNTO 22) WHEN x"00000016",
	"00000000000000000000000" & SrcA(31 DOWNTO 23) WHEN x"00000017",
	"000000000000000000000000" & SrcA(31 DOWNTO 24) WHEN x"00000018",
	"0000000000000000000000000" & SrcA(31 DOWNTO 25) WHEN x"00000019",
	"00000000000000000000000000" & SrcA(31 DOWNTO 26) WHEN x"0000001A",
	"000000000000000000000000000" & SrcA(31 DOWNTO 27) WHEN x"0000001B",
	"0000000000000000000000000000" & SrcA(31 DOWNTO 28) WHEN x"0000001C",
	"00000000000000000000000000000" & SrcA(31 DOWNTO 29) WHEN x"0000001D",
	"000000000000000000000000000000" & SrcA(31 DOWNTO 30) WHEN x"0000001E",
	"0000000000000000000000000000000" & SrcA(31) WHEN x"0000001F",
	x"00000000" WHEN OTHERS;
-------------------------------------
with ALUControl select--ALUControl signal comes from the CU depending on the current instruction
ALUResult <= 	SrcA+SrcB when "000",
					SrcA-SrcB when "001",
					SrcA and SrcB when "010",
					SrcA or SrcB when "011",
					SrcA nor SrcB when "100",
					shiftleft when "101",
					shiftright when "110",
					SrcA+SrcB when others;	

with z select
Zero <= 	'1' when x"00000000",
			'0' when others;	
with z(31) select
LessThan <= 	'1' when '1',
					'0' when others;
with z select					
GreatThan <= 	'0' when x"00000000",
					--not z(31) when others;
					'1' when others;
----------------------------
end Behavioral;

